module testemaquinas();


